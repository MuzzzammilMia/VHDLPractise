--Aim of the project is just go over a simple project in VHDL
-- To cover VHDL again
-- Link https://www.nandland.com/vhdl/tutorials/tutorial-modelsim-simulation-walkthrough.html

library ieee;
use ieee.std_logic_1164.all;
 
entity and_gate is
  port (
    input_1    : in  std_logic;
    input_2    : in  std_logic;
    and_result : out std_logic
    );
end and_gate;
 
architecture rtl of and_gate is
  signal and_gate : std_logic;
begin
  and_gate   <= input_1 and input_2;
  and_result <= and_gate;
end rtl ;
